
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mStateMachine is
end mStateMachine;

architecture Behavioral of mStateMachine is

begin


end Behavioral;

